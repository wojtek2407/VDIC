
module orange (input wire A, output wire B);
	
	assign B = ~A;
	
endmodule

