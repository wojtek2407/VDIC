
module orange_tb;
	
	wire A;
	wire B;

	orange u_orange (
		.A(A),
		.B(B)
		);
	
endmodule